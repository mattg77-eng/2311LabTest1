
module Lab3(
    input  [9:0] SW,       
    output [6:0] HEX5, HEX3, HEX1, HEX0 
);

    wire [3:0] A = SW[3:0];    
    wire [3:0] B = SW[7:4];     
    wire S = SW[8];             

    wire [3:0] B_mod;
    wire [3:0] SUM;
    wire cout;

    assign B_mod = B ^ {4{S}};  


    wire [3:0] carry;
    full_adder FA0 (A[0], B_mod[0], S, SUM[0], carry[0]);
    full_adder FA1 (A[1], B_mod[1], carry[0], SUM[1], carry[1]);
    full_adder FA2 (A[2], B_mod[2], carry[1], SUM[2], carry[2]);
    full_adder FA3 (A[3], B_mod[3], carry[2], SUM[3], carry[3]);
    assign cout = carry[3];


    reg [3:0] display_result;
    reg [6:0] HEX1_reg;

    always @(*) begin
        HEX1_reg = 7'b111_1111; 
        display_result = SUM;

        if (S == 0) begin
           if (cout == 1) HEX1_reg = 7'b111_1001; 
        end 
        else begin
        
            if (cout == 0) begin
                HEX1_reg = 7'b011_1111; 
                display_result = (~SUM + 1'b1); 
            end
        end
    end

    hex_decoder hexA (A, HEX5);
    hex_decoder hexB (B, HEX3);
    hex_decoder hexRes (display_result, HEX0);

    assign HEX1 = HEX1_reg;

endmodule


module full_adder(
    input a, b, cin,
    output sum, cout
);
    assign sum = a ^ b ^ cin;
    assign cout = (a & b) | (b & cin) | (a & cin);
endmodule


module hex_decoder(
    input [3:0] hex,
    output reg [6:0] seg
);
    always @(*) begin
        case (hex)
            4'h0: seg = 7'b100_0000;
            4'h1: seg = 7'b111_1001;
            4'h2: seg = 7'b010_0100;
            4'h3: seg = 7'b011_0000;
            4'h4: seg = 7'b001_1001;
            4'h5: seg = 7'b001_0010;
            4'h6: seg = 7'b000_0010;
            4'h7: seg = 7'b111_1000;
            4'h8: seg = 7'b000_0000;
            4'h9: seg = 7'b001_0000;
            4'hA: seg = 7'b000_1000;
            4'hB: seg = 7'b000_0011;
            4'hC: seg = 7'b100_0110;
            4'hD: seg = 7'b010_0001;
            4'hE: seg = 7'b000_0110;
            4'hF: seg = 7'b000_1110;
            default: seg = 7'b111_1111;
        endcase
    end
endmodule
